localparam SBUS_IMM      = 5'b00000,     //immediate
           SBUS_COMP_IMM = 5'b00001,	   //complement of immediate
	        SBUS_S_LOG    = 5'b00010,     //scalar logical
	        SBUS_S_SHIFT  = 5'b00011,     //scalar shift 
	        SBUS_S_ADD    = 5'b00100,     //scalar add
	        SBUS_FP_ADD   = 5'b00101,     //floating point add
	        SBUS_FP_MULT  = 5'b00110,     //floating point multiply
	        SBUS_FP_RA    = 5'b00111,     //floating point reciprocal approximation
	        SBUS_CONST_GEN= 5'b01000,     //transmit (Ak) or constant to Si
	        SBUS_RTC      = 5'b01001,     //real time clock
	        SBUS_V_MASK   = 5'b01010,     //vector mask
	        SBUS_T_BUS    = 5'b01011,     //transmit (Tjk) to Si
	        SBUS_V0       = 5'b01100,     //transmit (Vj) to Si
			  SBUS_V1       = 5'b01101,
			  SBUS_V2       = 5'b01110,
			  SBUS_V3       = 5'b01111,
			  SBUS_V4       = 5'b10000,
			  SBUS_V5       = 5'b10001,
			  SBUS_V6       = 5'b10010,
			  SBUS_V7       = 5'b10011,
	        SBUS_MEM      = 5'b10100,
   	     SBUS_NONE     = 5'b10101;
			  
			  
localparam ABUS_IMM      = 4'b0000,     //immediate
           ABUS_COMP_IMM = 4'b0001,	   //complement of immediate
	        ABUS_SIMM     = 4'b0010,     //short immediate
	        ABUS_S_BUS    = 4'b0011,     //transmit (Sj) to Ai
	        ABUS_B_BUS    = 4'b0100,     //transmit (Bjk) to Ai
	        ABUS_S_POP    = 4'b0101,     //scalar population count
	        ABUS_A_ADD    = 4'b0110,     //address add
	        ABUS_A_MULT   = 4'b0111,     //address multiply
	        ABUS_A_BUS    = 4'b1000,     //transmit (Ak) to Si
	        ABUS_CHANNEL  = 4'b1001,     //real time clock
	        ABUS_MEM      = 4'b1010,     //memory
   	     ABUS_NONE     = 4'b1011;
